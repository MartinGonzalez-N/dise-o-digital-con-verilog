module soluciones (input IN_A, IN_B, IN_C, IN_D, output a, b, c, d, e, f, g);
	display dis(.num_0(IN_A),.num_1(IN_B),.num_2(IN_C),.num_3(IN_D),.a(a),.b(b),.c(c),.d(d),.e(e),.f(f),.g(g));
endmodule
